** Profile: "SCHEMATIC1-orcad8week4"  [ C:\Users\OHSEHOON\Desktop\pispice\orcad8week4-PSpiceFiles\SCHEMATIC1\orcad8week4.sim ] 

** Creating circuit file "orcad8week4.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\OHSEHOON\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 2m 0 
.STEP PARAM cval LIST 0.001u, 0.01u, 0.1u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
