** Profile: "SCHEMATIC1-orcad13week11"  [ C:\Users\OHSEHOON\Desktop\pispice\orcad13week11-PSpiceFiles\SCHEMATIC1\orcad13week11.sim ] 

** Creating circuit file "orcad13week11.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "C:\Users\OHSEHOON\Desktop\pispice\orcad13week11-PSpiceFiles\SCHEMATIC1\orcad13week11\orcad13week11_profile.inc" 
* Local Libraries :
.STMLIB "../../../orcad13week11-pspicefiles/orcad13week11.stl" 
* From [PSPICE NETLIST] section of C:\Users\OHSEHOON\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
