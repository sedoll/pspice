** Profile: "SCHEMATIC1-orcad13week4"  [ C:\Users\OHSEHOON\Desktop\pispice\orcad13week4-PSpiceFiles\SCHEMATIC1\orcad13week4.sim ] 

** Creating circuit file "orcad13week4.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "../../../orcad13week4-PSpiceFiles/ORCAD13WEEK4.stl" 
* From [PSPICE NETLIST] section of C:\Users\OHSEHOON\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1200ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
