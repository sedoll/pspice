** Profile: "SCHEMATIC1-orcad7week1"  [ C:\Users\OHSEHOON\Desktop\pispice\orcad7week1-PSpiceFiles\SCHEMATIC1\orcad7week1.sim ] 

** Creating circuit file "orcad7week1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../orcad7week1-pspicefiles/orcad7week1.lib" 
* From [PSPICE NETLIST] section of C:\Users\OHSEHOON\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN PARAM P 0 5 0.1 
.MC 10 DC I(V_Meter) YMAX OUTPUT ALL 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
