** Profile: "SCHEMATIC1-orcad13week10"  [ C:\Users\OHSEHOON\Desktop\pispice\orcad13week10-PSpiceFiles\SCHEMATIC1\orcad13week10.sim ] 

** Creating circuit file "orcad13week10.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "../../../orcad13week10-PSpiceFiles/ORCAD13WEEK10.stl" 
* From [PSPICE NETLIST] section of C:\Users\OHSEHOON\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1.6u 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
