** Profile: "SCHEMATIC1-orcad14week6"  [ C:\Users\OHSEHOON\Desktop\pispice\orcad14week6-PSpiceFiles\SCHEMATIC1\orcad14week6.sim ] 

** Creating circuit file "orcad14week6.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\OHSEHOON\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V5 0 -10 -1 
.STEP LIN V_V6 -3.5 -5 -0.5 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
