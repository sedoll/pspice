** Profile: "SCHEMATIC1-orcad8week2"  [ C:\Users\OHSEHOON\Desktop\pispice\orcad8week2-PSpiceFiles\SCHEMATIC1\orcad8week2.sim ] 

** Creating circuit file "orcad8week2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\OHSEHOON\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 2.5m 0 
.STEP PARAM rval LIST 1k, 10k, 100k 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
