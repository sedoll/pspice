** Profile: "SCHEMATIC1-orcad10week5"  [ C:\Users\OHSEHOON\Desktop\pispice\orcad10week5-PSpiceFiles\SCHEMATIC1\orcad10week5.sim ] 

** Creating circuit file "orcad10week5.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\OHSEHOON\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V1 -1 0.5 0.01 
.STEP TEMP LIST -10, 0, 10 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
