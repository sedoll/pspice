** Profile: "SCHEMATIC1-orcad13week5"  [ C:\Users\OHSEHOON\Desktop\pispice\orcad13week6-PSpiceFiles\SCHEMATIC1\orcad13week5.sim ] 

** Creating circuit file "orcad13week5.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "../../../orcad13week6-PSpiceFiles/ORCAD13WEEK6.stl" 
* From [PSPICE NETLIST] section of C:\Users\OHSEHOON\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
