** Profile: "SCHEMATIC1-orcad10week4"  [ C:\Users\OHSEHOON\Desktop\pispice\orcad10week4-PSpiceFiles\SCHEMATIC1\orcad10week4.sim ] 

** Creating circuit file "orcad10week4.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\OHSEHOON\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V1 -1 2 0.01 
.STEP TEMP LIST -100, 0, 100 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
